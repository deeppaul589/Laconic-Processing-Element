`timescale 1ns / 1ps

module tb();
    
    reg [15:0] in_applied;
    reg [47:0] t0;
    reg [47:0] t1;
    reg [15:0] s0;
    reg [15:0] s1;
    
    wire signed [21:0] result;
    
    core uut(
    
        .in_applied(in_applied),
        .t0(t0),
        .t1(t1),
        .s0(s0),
        .s1(s1),
        .out_value(result)
    
    );
    
    
    
    initial begin
        
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd0, 3'd2, 3'd7, 3'd0, 3'd2, 3'd7, 3'd0, 3'd2, 3'd7, 3'd0, 3'd2, 3'd5, 3'd7, 3'd0, 3'd2, 3'd5};
t1 = {3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd4, 3'd4, 3'd4, 3'd3, 3'd3, 3'd3, 3'd3, 3'd7, 3'd7, 3'd7};
s0 = {1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0};
s1 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1};
//MAC result =  -1889
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd7, 3'd1, 3'd3, 3'd5, 3'd1, 3'd3, 3'd5, 3'd1, 3'd3, 3'd5, 3'd0, 3'd1, 3'd6, 3'd0, 3'd1, 3'd6};
t1 = {3'd7, 3'd0, 3'd0, 3'd0, 3'd2, 3'd2, 3'd2, 3'd6, 3'd6, 3'd6, 3'd0, 3'd0, 3'd0, 3'd4, 3'd4, 3'd4};
s0 = {1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
s1 = {1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
//MAC result =  20085
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd0, 3'd1, 3'd6, 3'd1, 3'd3, 3'd5, 3'd1, 3'd3, 3'd5, 3'd1, 3'd3, 3'd5, 3'd0, 3'd3, 3'd5, 3'd6};
t1 = {3'd6, 3'd6, 3'd6, 3'd0, 3'd0, 3'd0, 3'd2, 3'd2, 3'd2, 3'd6, 3'd6, 3'd6, 3'd0, 3'd0, 3'd0, 3'd0};
s0 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1};
s1 = {1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0};
//MAC result =  -7191
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd0, 3'd3, 3'd5, 3'd6, 3'd0, 3'd3, 3'd5, 3'd6, 3'd4, 3'd7, 3'd4, 3'd7, 3'd0, 3'd5, 3'd0, 3'd5};
t1 = {3'd3, 3'd3, 3'd3, 3'd3, 3'd6, 3'd6, 3'd6, 3'd6, 3'd2, 3'd2, 3'd6, 3'd6, 3'd0, 3'd0, 3'd5, 3'd5};
s0 = {1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b0};
s1 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0};
//MAC result =  2201
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd0, 3'd2, 3'd5, 3'd7, 3'd0, 3'd4, 3'd7, 3'd0, 3'd4, 3'd7, 3'd0, 3'd4, 3'd7, 3'd1, 3'd5, 3'd1};
t1 = {3'd6, 3'd6, 3'd6, 3'd6, 3'd2, 3'd2, 3'd2, 3'd4, 3'd4, 3'd4, 3'd7, 3'd7, 3'd7, 3'd1, 3'd1, 3'd4};
s0 = {1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1};
s1 = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1};
//MAC result =  18296
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd5, 3'd0, 3'd3, 3'd4, 3'd6, 3'd0, 3'd3, 3'd4, 3'd6, 3'd2, 3'd3, 3'd7, 3'd2, 3'd3, 3'd7, 3'd2};
t1 = {3'd4, 3'd1, 3'd1, 3'd1, 3'd1, 3'd6, 3'd6, 3'd6, 3'd6, 3'd3, 3'd3, 3'd3, 3'd5, 3'd5, 3'd5, 3'd6};
s0 = {1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0};
s1 = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1};
//MAC result =  -142
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd3, 3'd7, 3'd5, 3'd6, 3'd5, 3'd6, 3'd5, 3'd6, 3'd1, 3'd2, 3'd5, 3'd6, 3'd1, 3'd2, 3'd5, 3'd6};
t1 = {3'd6, 3'd6, 3'd0, 3'd0, 3'd5, 3'd5, 3'd7, 3'd7, 3'd4, 3'd4, 3'd4, 3'd4, 3'd6, 3'd6, 3'd6, 3'd6};
s0 = {1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
s1 = {1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1};
//MAC result =  -6528
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0};
t0 = {3'd1, 3'd3, 3'd7, 3'd1, 3'd3, 3'd7, 3'd1, 3'd3, 3'd7, 3'd0, 3'd5, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0};
t1 = {3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd4, 3'd4, 3'd4, 3'd0, 3'd0, 3'd5, 3'd5, 3'd0, 3'd0, 3'd0};
s0 = {1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1};
s1 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1};
//MAC result =  -1281
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd0, 3'd3, 3'd4, 3'd6, 3'd0, 3'd3, 3'd4, 3'd6, 3'd2, 3'd2, 3'd0, 3'd4, 3'd6, 3'd0, 3'd4, 3'd6};
t1 = {3'd2, 3'd2, 3'd2, 3'd2, 3'd6, 3'd6, 3'd6, 3'd6, 3'd0, 3'd4, 3'd0, 3'd0, 3'd0, 3'd2, 3'd2, 3'd2};
s0 = {1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0};
s1 = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
//MAC result =  -5461
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd0, 3'd4, 3'd6, 3'd0, 3'd4, 3'd6, 3'd3, 3'd4, 3'd6, 3'd0, 3'd2, 3'd6, 3'd0, 3'd2, 3'd6, 3'd0};
t1 = {3'd4, 3'd4, 3'd4, 3'd7, 3'd7, 3'd7, 3'd3, 3'd3, 3'd3, 3'd2, 3'd2, 3'd2, 3'd4, 3'd4, 3'd4, 3'd7};
s0 = {1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
s1 = {1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0};
//MAC result =  10804
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd2, 3'd6, 3'd0, 3'd2, 3'd7, 3'd0, 3'd2, 3'd7, 3'd0, 3'd2, 3'd7, 3'd2, 3'd4, 3'd6, 3'd2, 3'd4};
t1 = {3'd7, 3'd7, 3'd0, 3'd0, 3'd0, 3'd2, 3'd2, 3'd2, 3'd6, 3'd6, 3'd6, 3'd2, 3'd2, 3'd2, 3'd5, 3'd5};
s0 = {1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0};
s1 = {1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0};
//MAC result =  375
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0};
t0 = {3'd6, 3'd2, 3'd4, 3'd6, 3'd2, 3'd5, 3'd2, 3'd5, 3'd0, 3'd5, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0};
t1 = {3'd5, 3'd6, 3'd6, 3'd6, 3'd4, 3'd4, 3'd6, 3'd6, 3'd0, 3'd0, 3'd5, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0};
s0 = {1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1};
s1 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1};
//MAC result =  -5727
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd2, 3'd5, 3'd6, 3'd2, 3'd5, 3'd6, 3'd2, 3'd5, 3'd6, 3'd2, 3'd5, 3'd6, 3'd2, 3'd6, 3'd2, 3'd6};
t1 = {3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd5, 3'd5, 3'd5, 3'd7, 3'd7, 3'd7, 3'd0, 3'd0, 3'd5, 3'd5};
s0 = {1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
s1 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0};
//MAC result =  1368
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd2, 3'd6, 3'd0, 3'd5, 3'd0, 3'd5, 3'd0, 3'd5, 3'd0, 3'd5, 3'd0, 3'd2, 3'd5, 3'd6, 3'd0, 3'd2};
t1 = {3'd6, 3'd6, 3'd1, 3'd1, 3'd4, 3'd4, 3'd5, 3'd5, 3'd7, 3'd7, 3'd2, 3'd2, 3'd2, 3'd2, 3'd3, 3'd3};
s0 = {1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1};
s1 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
//MAC result =  -6934
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd5, 3'd6, 3'd0, 3'd2, 3'd5, 3'd6, 3'd0, 3'd5, 3'd6, 3'd0, 3'd5, 3'd6, 3'd0, 3'd5, 3'd6, 3'd0};
t1 = {3'd3, 3'd3, 3'd7, 3'd7, 3'd7, 3'd7, 3'd2, 3'd2, 3'd2, 3'd4, 3'd4, 3'd4, 3'd6, 3'd6, 3'd6, 3'd1};
s0 = {1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b0};
s1 = {1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1};
//MAC result =  5674
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd2, 3'd7, 3'd0, 3'd2, 3'd7, 3'd0, 3'd2, 3'd7, 3'd2, 3'd4, 3'd7, 3'd2, 3'd4, 3'd7, 3'd1, 3'd4};
t1 = {3'd1, 3'd1, 3'd4, 3'd4, 3'd4, 3'd6, 3'd6, 3'd6, 3'd4, 3'd4, 3'd4, 3'd5, 3'd5, 3'd5, 3'd0, 3'd0};
s0 = {1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0};
s1 = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1};
//MAC result =  -4694
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0};
t0 = {3'd6, 3'd1, 3'd4, 3'd6, 3'd1, 3'd4, 3'd6, 3'd1, 3'd4, 3'd6, 3'd0, 3'd5, 3'd0, 3'd5, 3'd0, 3'd0};
t1 = {3'd0, 3'd3, 3'd3, 3'd3, 3'd4, 3'd4, 3'd4, 3'd7, 3'd7, 3'd7, 3'd0, 3'd0, 3'd5, 3'd5, 3'd0, 3'd0};
s0 = {1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1};
s1 = {1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1};
//MAC result =  -4943
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd1, 3'd3, 3'd4, 3'd1, 3'd3, 3'd4, 3'd1, 3'd3, 3'd4, 3'd0, 3'd5, 3'd6, 3'd0, 3'd5, 3'd6, 3'd0};
t1 = {3'd0, 3'd0, 3'd0, 3'd3, 3'd3, 3'd3, 3'd5, 3'd5, 3'd5, 3'd0, 3'd0, 3'd0, 3'd2, 3'd2, 3'd2, 3'd5};
s0 = {1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1};
s1 = {1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
//MAC result =  53
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd5, 3'd6, 3'd3, 3'd6, 3'd7, 3'd3, 3'd6, 3'd7, 3'd3, 3'd6, 3'd7, 3'd3, 3'd6, 3'd7, 3'd0, 3'd3};
t1 = {3'd5, 3'd5, 3'd0, 3'd0, 3'd0, 3'd2, 3'd2, 3'd2, 3'd3, 3'd3, 3'd3, 3'd7, 3'd7, 3'd7, 3'd4, 3'd4};
s0 = {1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0};

s1 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
//MAC result =  5272
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd5, 3'd7, 3'd0, 3'd3, 3'd5, 3'd7, 3'd0, 3'd2, 3'd5, 3'd7, 3'd0, 3'd2, 3'd5, 3'd7, 3'd1, 3'd4};
t1 = {3'd4, 3'd4, 3'd7, 3'd7, 3'd7, 3'd7, 3'd2, 3'd2, 3'd2, 3'd2, 3'd4, 3'd4, 3'd4, 3'd4, 3'd1, 3'd1};
s0 = {1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0};
s1 = {1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
//MAC result =  -11520
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd1, 3'd4, 3'd0, 3'd3, 3'd6, 3'd7, 3'd0, 3'd3, 3'd6, 3'd7, 3'd0, 3'd3, 3'd6, 3'd7, 3'd0, 3'd5};
t1 = {3'd7, 3'd7, 3'd1, 3'd1, 3'd1, 3'd1, 3'd2, 3'd2, 3'd2, 3'd2, 3'd4, 3'd4, 3'd4, 3'd4, 3'd0, 3'd0};
s0 = {1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0};
s1 = {1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1};
//MAC result =  -3033
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
t0 = {3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0};
t1 = {3'd5, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0};
s0 = {1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
s1 = {1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
//MAC result =  992
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd2, 3'd4, 3'd5, 3'd0, 3'd3, 3'd4, 3'd6, 3'd0, 3'd3, 3'd4, 3'd6, 3'd0, 3'd3, 3'd4, 3'd6, 3'd0};
t1 = {3'd5, 3'd5, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd2, 3'd2, 3'd2, 3'd5, 3'd5, 3'd5, 3'd5, 3'd7};
s0 = {1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1};
s1 = {1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1};
//MAC result =  -2725
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd3, 3'd4, 3'd6, 3'd1, 3'd4, 3'd6, 3'd7, 3'd2, 3'd6, 3'd2, 3'd6, 3'd2, 3'd6, 3'd1, 3'd5, 3'd7};
t1 = {3'd7, 3'd7, 3'd7, 3'd2, 3'd2, 3'd2, 3'd2, 3'd0, 3'd0, 3'd4, 3'd4, 3'd6, 3'd6, 3'd0, 3'd0, 3'd0};
s0 = {1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1};
s1 = {1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0};
//MAC result =  98
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd1, 3'd5, 3'd7, 3'd1, 3'd5, 3'd7, 3'd0, 3'd1, 3'd5, 3'd6, 3'd0, 3'd1, 3'd5, 3'd6, 3'd0, 3'd1};
t1 = {3'd2, 3'd2, 3'd2, 3'd7, 3'd7, 3'd7, 3'd0, 3'd0, 3'd0, 3'd0, 3'd3, 3'd3, 3'd3, 3'd3, 3'd6, 3'd6};
s0 = {1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
s1 = {1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
//MAC result =  13235
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd5, 3'd6, 3'd0, 3'd1, 3'd5, 3'd6, 3'd0, 3'd1, 3'd6, 3'd0, 3'd1, 3'd6, 3'd0, 3'd1, 3'd6, 3'd3};
t1 = {3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd1, 3'd1, 3'd1, 3'd2, 3'd2, 3'd2, 3'd6, 3'd6, 3'd6, 3'd0};
s0 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
s1 = {1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0};
//MAC result =  -11210
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0};
t0 = {3'd4, 3'd7, 3'd3, 3'd4, 3'd7, 3'd3, 3'd4, 3'd7, 3'd0, 3'd5, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0};
t1 = {3'd0, 3'd0, 3'd2, 3'd2, 3'd2, 3'd5, 3'd5, 3'd5, 3'd0, 3'd0, 3'd5, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0};
s0 = {1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1};
s1 = {1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1};
//MAC result =  -2031
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd4, 3'd7, 3'd4, 3'd7, 3'd2, 3'd5, 3'd6, 3'd2, 3'd5, 3'd6, 3'd2, 3'd5, 3'd6, 3'd1, 3'd5, 3'd6};
t1 = {3'd2, 3'd2, 3'd5, 3'd5, 3'd1, 3'd1, 3'd1, 3'd4, 3'd4, 3'd4, 3'd6, 3'd6, 3'd6, 3'd0, 3'd0, 3'd0};
s0 = {1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0};
s1 = {1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
//MAC result =  11942
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd1, 3'd5, 3'd6, 3'd1, 3'd5, 3'd6, 3'd3, 3'd3, 3'd2, 3'd2, 3'd4, 3'd6, 3'd4, 3'd6, 3'd4, 3'd6};
t1 = {3'd4, 3'd4, 3'd4, 3'd6, 3'd6, 3'd6, 3'd3, 3'd7, 3'd0, 3'd6, 3'd0, 3'd0, 3'd3, 3'd3, 3'd4, 3'd4};
s0 = {1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1};
s1 = {1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1};
//MAC result =  -2188
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd1, 3'd4, 3'd6, 3'd1, 3'd4, 3'd6, 3'd1, 3'd4, 3'd6, 3'd1, 3'd2, 3'd5, 3'd7, 3'd1, 3'd2, 3'd5};
t1 = {3'd1, 3'd1, 3'd1, 3'd3, 3'd3, 3'd3, 3'd4, 3'd4, 3'd4, 3'd2, 3'd2, 3'd2, 3'd2, 3'd4, 3'd4, 3'd4};
s0 = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0};
s1 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
//MAC result =  -2380
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
t0 = {3'd7, 3'd0, 3'd5, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0};
t1 = {3'd4, 3'd0, 3'd0, 3'd5, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0};
s0 = {1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
s1 = {1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
//MAC result =  3009
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd0, 3'd0, 3'd0, 3'd0, 3'd3, 3'd5, 3'd6, 3'd0, 3'd3, 3'd5, 3'd6, 3'd1, 3'd2, 3'd4, 3'd7, 3'd1};
t1 = {3'd0, 3'd3, 3'd6, 3'd0, 3'd0, 3'd0, 3'd0, 3'd5, 3'd5, 3'd5, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd3};
s0 = {1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0};
s1 = {1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0};
//MAC result =  -2564
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd2, 3'd4, 3'd7, 3'd1, 3'd2, 3'd4, 3'd7, 3'd1, 3'd2, 3'd4, 3'd7, 3'd0, 3'd1, 3'd4, 3'd6, 3'd0};
t1 = {3'd3, 3'd3, 3'd3, 3'd5, 3'd5, 3'd5, 3'd5, 3'd6, 3'd6, 3'd6, 3'd6, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2};
s0 = {1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
s1 = {1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1};
//MAC result =  9391
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd1, 3'd4, 3'd6, 3'd0, 3'd1, 3'd4, 3'd6, 3'd0, 3'd1, 3'd4, 3'd6, 3'd3, 3'd5, 3'd7, 3'd3, 3'd5};
t1 = {3'd2, 3'd2, 3'd2, 3'd4, 3'd4, 3'd4, 3'd4, 3'd6, 3'd6, 3'd6, 3'd6, 3'd0, 3'd0, 3'd0, 3'd4, 3'd4};
s0 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0};
s1 = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
//MAC result =  -6416
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd7, 3'd3, 3'd5, 3'd7, 3'd4, 3'd6, 3'd2, 3'd2, 3'd2, 3'd1, 3'd5, 3'd6, 3'd1, 3'd5, 3'd6, 3'd0};
t1 = {3'd4, 3'd6, 3'd6, 3'd6, 3'd4, 3'd4, 3'd0, 3'd2, 3'd4, 3'd2, 3'd2, 3'd2, 3'd4, 3'd4, 3'd4, 3'd0};
s0 = {1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1};
s1 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1};
//MAC result =  -9587
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
t0 = {3'd5, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0};
t1 = {3'd0, 3'd5, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0};
s0 = {1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
s1 = {1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
//MAC result =  992
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd0, 3'd2, 3'd4, 3'd6, 3'd0, 3'd2, 3'd4, 3'd6, 3'd0, 3'd2, 3'd4, 3'd6, 3'd2, 3'd6, 3'd2, 3'd6};
t1 = {3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd4, 3'd4, 3'd4, 3'd6, 3'd6, 3'd6, 3'd6, 3'd1, 3'd1, 3'd4, 3'd4};
s0 = {1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b0};
s1 = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1};
//MAC result =  -4981
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd2, 3'd6, 3'd0, 3'd3, 3'd4, 3'd6, 3'd1, 3'd0, 3'd4, 3'd0, 3'd4, 3'd0, 3'd4, 3'd0, 3'd4, 3'd2};
t1 = {3'd6, 3'd6, 3'd0, 3'd0, 3'd0, 3'd0, 3'd7, 3'd0, 3'd0, 3'd2, 3'd2, 3'd4, 3'd4, 3'd6, 3'd6, 3'd2};
s0 = {1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
s1 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0};
//MAC result =  5476
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd5, 3'd7, 3'd2, 3'd5, 3'd7, 3'd0, 3'd2, 3'd4, 3'd7, 3'd0, 3'd2, 3'd4, 3'd7, 3'd0, 3'd2, 3'd4};
t1 = {3'd2, 3'd2, 3'd6, 3'd6, 3'd6, 3'd1, 3'd1, 3'd1, 3'd1, 3'd4, 3'd4, 3'd4, 3'd4, 3'd5, 3'd5, 3'd5};
s0 = {1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1};

s1 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
//MAC result =  -5130
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0};
t0 = {3'd7, 3'd0, 3'd2, 3'd4, 3'd7, 3'd2, 3'd3, 3'd5, 3'd2, 3'd3, 3'd5, 3'd0, 3'd5, 3'd0, 3'd5, 3'd0};
t1 = {3'd5, 3'd6, 3'd6, 3'd6, 3'd6, 3'd4, 3'd4, 3'd4, 3'd6, 3'd6, 3'd6, 3'd0, 3'd0, 3'd5, 3'd5, 3'd0};
s0 = {1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1};
s1 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1};
//MAC result =  15937
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd2, 3'd4, 3'd6, 3'd2, 3'd4, 3'd6, 3'd2, 3'd4, 3'd6, 3'd0, 3'd3, 3'd6, 3'd0, 3'd3, 3'd6, 3'd0};
t1 = {3'd0, 3'd0, 3'd0, 3'd2, 3'd2, 3'd2, 3'd4, 3'd4, 3'd4, 3'd2, 3'd2, 3'd2, 3'd4, 3'd4, 3'd4, 3'd5};
s0 = {1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
s1 = {1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
//MAC result =  2480
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd3, 3'd6, 3'd0, 3'd2, 3'd6, 3'd0, 3'd2, 3'd6, 3'd0, 3'd2, 3'd6, 3'd0, 3'd2, 3'd6, 3'd0, 3'd2};
t1 = {3'd5, 3'd5, 3'd1, 3'd1, 3'd1, 3'd2, 3'd2, 3'd2, 3'd4, 3'd4, 3'd4, 3'd7, 3'd7, 3'd7, 3'd1, 3'd1};
s0 = {1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0};
s1 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
//MAC result =  8760
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd7, 3'd0, 3'd2, 3'd7, 3'd1, 3'd2, 3'd4, 3'd1, 3'd2, 3'd4, 3'd5, 3'd6, 3'd5, 3'd6, 3'd1, 3'd4};
t1 = {3'd1, 3'd6, 3'd6, 3'd6, 3'd1, 3'd1, 3'd1, 3'd5, 3'd5, 3'd5, 3'd1, 3'd1, 3'd6, 3'd6, 3'd4, 3'd4};
s0 = {1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
s1 = {1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1};
//MAC result =  14540
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0};
t0 = {3'd6, 3'd7, 3'd2, 3'd7, 3'd2, 3'd7, 3'd2, 3'd7, 3'd0, 3'd5, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0};
t1 = {3'd4, 3'd4, 3'd1, 3'd1, 3'd2, 3'd2, 3'd4, 3'd4, 3'd0, 3'd0, 3'd5, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0};
s0 = {1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1};
s1 = {1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1};
//MAC result =  281
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd1, 3'd2, 3'd5, 3'd7, 3'd2, 3'd4, 3'd2, 3'd4, 3'd0, 3'd5, 3'd6, 3'd0, 3'd5, 3'd6, 3'd0, 3'd5};
t1 = {3'd4, 3'd4, 3'd4, 3'd4, 3'd1, 3'd1, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd4, 3'd4, 3'd4, 3'd6, 3'd6};
s0 = {1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0};
s1 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
//MAC result =  -2908
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd6, 3'd1, 3'd2, 3'd1, 3'd2, 3'd1, 3'd2, 3'd1, 3'd2, 3'd1, 3'd4, 3'd7, 3'd1, 3'd4, 3'd7, 3'd1};
t1 = {3'd6, 3'd0, 3'd0, 3'd3, 3'd3, 3'd4, 3'd4, 3'd6, 3'd6, 3'd1, 3'd1, 3'd1, 3'd2, 3'd2, 3'd2, 3'd5};
s0 = {1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0};
s1 = {1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
//MAC result =  3958
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd4, 3'd7, 3'd1, 3'd4, 3'd6, 3'd1, 3'd4, 3'd6, 3'd1, 3'd4, 3'd6, 3'd0, 3'd1, 3'd4, 3'd0, 3'd1};
t1 = {3'd5, 3'd5, 3'd2, 3'd2, 3'd2, 3'd5, 3'd5, 3'd5, 3'd6, 3'd6, 3'd6, 3'd1, 3'd1, 3'd1, 3'd5, 3'd5};
s0 = {1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
s1 = {1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0};
//MAC result =  -8126
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0};
t0 = {3'd4, 3'd0, 3'd1, 3'd4, 3'd4, 3'd7, 3'd4, 3'd7, 3'd0, 3'd5, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0};
t1 = {3'd5, 3'd6, 3'd6, 3'd6, 3'd0, 3'd0, 3'd6, 3'd6, 3'd0, 3'd0, 3'd5, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0};
s0 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1};
s1 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1};
//MAC result =  -4335
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd0, 3'd2, 3'd4, 3'd7, 3'd0, 3'd2, 3'd4, 3'd7, 3'd0, 3'd2, 3'd4, 3'd7, 3'd4, 3'd4, 3'd3, 3'd5};
t1 = {3'd0, 3'd0, 3'd0, 3'd0, 3'd3, 3'd3, 3'd3, 3'd3, 3'd4, 3'd4, 3'd4, 3'd4, 3'd0, 3'd3, 3'd0, 3'd0};
s0 = {1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0};
s1 = {1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0};
//MAC result =  -2309
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd3, 3'd5, 3'd3, 3'd5, 3'd3, 3'd5, 3'd3, 3'd6, 3'd3, 3'd6, 3'd3, 3'd6, 3'd0, 3'd5, 3'd7, 3'd0};
t1 = {3'd3, 3'd3, 3'd4, 3'd4, 3'd6, 3'd6, 3'd1, 3'd1, 3'd2, 3'd2, 3'd7, 3'd7, 3'd0, 3'd0, 3'd0, 3'd1};
s0 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0};
s1 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0};
//MAC result =  11699
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd5, 3'd7, 3'd0, 3'd5, 3'd7, 3'd0, 3'd5, 3'd7, 3'd2, 3'd4, 3'd6, 3'd2, 3'd4, 3'd6, 3'd1, 3'd4};
t1 = {3'd1, 3'd1, 3'd3, 3'd3, 3'd3, 3'd7, 3'd7, 3'd7, 3'd1, 3'd1, 3'd1, 3'd7, 3'd7, 3'd7, 3'd1, 3'd1};
s0 = {1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1};
s1 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
//MAC result =  16788
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0};
t0 = {3'd6, 3'd1, 3'd4, 3'd6, 3'd1, 3'd4, 3'd6, 3'd4, 3'd6, 3'd4, 3'd6, 3'd0, 3'd5, 3'd0, 3'd5, 3'd0};
t1 = {3'd1, 3'd4, 3'd4, 3'd4, 3'd6, 3'd6, 3'd6, 3'd1, 3'd1, 3'd3, 3'd3, 3'd0, 3'd0, 3'd5, 3'd5, 3'd0};
s0 = {1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1};
s1 = {1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1};
//MAC result =  -2175
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd4, 3'd6, 3'd4, 3'd6, 3'd5, 3'd7, 3'd5, 3'd7, 3'd5, 3'd7, 3'd1, 3'd4, 3'd6, 3'd1, 3'd4, 3'd6};
t1 = {3'd3, 3'd3, 3'd7, 3'd7, 3'd0, 3'd0, 3'd2, 3'd2, 3'd7, 3'd7, 3'd0, 3'd0, 3'd0, 3'd5, 3'd5, 3'd5};
s0 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0};
s1 = {1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
//MAC result =  -18834
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd1, 3'd4, 3'd6, 3'd0, 3'd5, 3'd0, 3'd5, 3'd0, 3'd5, 3'd0, 3'd5, 3'd0, 3'd7, 3'd0, 3'd7, 3'd0};
t1 = {3'd6, 3'd6, 3'd6, 3'd0, 3'd0, 3'd2, 3'd2, 3'd4, 3'd4, 3'd6, 3'd6, 3'd0, 3'd0, 3'd3, 3'd3, 3'd0};
s0 = {1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1};
s1 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1};
//MAC result =  7469
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd3, 3'd6, 3'd0, 3'd3, 3'd6, 3'd0, 3'd3, 3'd6, 3'd0, 3'd3, 3'd6, 3'd0, 3'd2, 3'd3, 3'd5, 3'd0};
t1 = {3'd0, 3'd0, 3'd2, 3'd2, 3'd2, 3'd4, 3'd4, 3'd4, 3'd6, 3'd6, 3'd6, 3'd2, 3'd2, 3'd2, 3'd2, 3'd6};
s0 = {1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
s1 = {1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1};
//MAC result =  4504
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
t0 = {3'd2, 3'd3, 3'd5, 3'd0, 3'd5, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0};
t1 = {3'd6, 3'd6, 3'd6, 3'd0, 3'd0, 3'd5, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0};
s0 = {1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
s1 = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
//MAC result =  -1855
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd1, 3'd2, 3'd7, 3'd1, 3'd2, 3'd7, 3'd0, 3'd1, 3'd3, 3'd7, 3'd0, 3'd1, 3'd3, 3'd7, 3'd0, 3'd1};
t1 = {3'd2, 3'd2, 3'd2, 3'd6, 3'd6, 3'd6, 3'd3, 3'd3, 3'd3, 3'd3, 3'd5, 3'd5, 3'd5, 3'd5, 3'd6, 3'd6};

s0 = {1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0};
s1 = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
//MAC result =  -12784
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd3, 3'd7, 3'd1, 3'd4, 3'd6, 3'd1, 3'd4, 3'd6, 3'd1, 3'd4, 3'd6, 3'd2, 3'd5, 3'd6, 3'd2, 3'd5};
t1 = {3'd6, 3'd6, 3'd2, 3'd2, 3'd2, 3'd5, 3'd5, 3'd5, 3'd6, 3'd6, 3'd6, 3'd0, 3'd0, 3'd0, 3'd4, 3'd4};
s0 = {1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0};
s1 = {1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0};
//MAC result =  -10148
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd6, 3'd2, 3'd5, 3'd6, 3'd0, 3'd1, 3'd2, 3'd5, 3'd0, 3'd1, 3'd2, 3'd5, 3'd0, 3'd1, 3'd2, 3'd5};
t1 = {3'd4, 3'd6, 3'd6, 3'd6, 3'd2, 3'd2, 3'd2, 3'd2, 3'd5, 3'd5, 3'd5, 3'd5, 3'd6, 3'd6, 3'd6, 3'd6};
s0 = {1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
s1 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1};
//MAC result =  -4732
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd4, 3'd7, 3'd4, 3'd7, 3'd4, 3'd7, 3'd4, 3'd7, 3'd0, 3'd3, 3'd5, 3'd6, 3'd0, 3'd3, 3'd5, 3'd6};
t1 = {3'd0, 3'd0, 3'd2, 3'd2, 3'd4, 3'd4, 3'd6, 3'd6, 3'd0, 3'd0, 3'd0, 3'd0, 3'd3, 3'd3, 3'd3, 3'd3};
s0 = {1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1};
s1 = {1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0};
//MAC result =  8351
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd0, 3'd3, 3'd5, 3'd6, 3'd0, 3'd3, 3'd5, 3'd6, 3'd5, 3'd7, 3'd5, 3'd7, 3'd5, 3'd7, 3'd5, 3'd7};
t1 = {3'd5, 3'd5, 3'd5, 3'd5, 3'd6, 3'd6, 3'd6, 3'd6, 3'd0, 3'd0, 3'd2, 3'd2, 3'd5, 3'd5, 3'd6, 3'd6};
s0 = {1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1};
s1 = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1};
//MAC result =  7296
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
t0 = {3'd0, 3'd5, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0};
t1 = {3'd0, 3'd0, 3'd5, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0};
s0 = {1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
s1 = {1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
//MAC result =  993
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd0, 3'd3, 3'd0, 3'd3, 3'd6, 3'd0, 3'd2, 3'd4, 3'd6, 3'd0, 3'd2, 3'd4, 3'd6, 3'd0, 3'd2, 3'd4};
t1 = {3'd1, 3'd1, 3'd5, 3'd5, 3'd5, 3'd3, 3'd3, 3'd3, 3'd3, 3'd5, 3'd5, 3'd5, 3'd5, 3'd6, 3'd6, 3'd6};
s0 = {1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0};
s1 = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
//MAC result =  838
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd6, 3'd0, 3'd3, 3'd4, 3'd0, 3'd3, 3'd4, 3'd0, 3'd3, 3'd4, 3'd1, 3'd3, 3'd5, 3'd1, 3'd3, 3'd5};
t1 = {3'd6, 3'd0, 3'd0, 3'd0, 3'd4, 3'd4, 3'd4, 3'd5, 3'd5, 3'd5, 3'd0, 3'd0, 3'd0, 3'd4, 3'd4, 3'd4};
s0 = {1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1};
s1 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0};
//MAC result =  -5613
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd1, 3'd3, 3'd5, 3'd0, 3'd2, 3'd3, 3'd6, 3'd0, 3'd2, 3'd6, 3'd0, 3'd2, 3'd6, 3'd0, 3'd2, 3'd6};
t1 = {3'd7, 3'd7, 3'd7, 3'd4, 3'd4, 3'd4, 3'd4, 3'd1, 3'd1, 3'd1, 3'd4, 3'd4, 3'd4, 3'd5, 3'd5, 3'd5};
s0 = {1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
s1 = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
//MAC result =  -1354
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd0, 3'd2, 3'd6, 3'd1, 3'd5, 3'd6, 3'd1, 3'd5, 3'd6, 3'd1, 3'd5, 3'd6, 3'd0, 3'd5, 3'd0, 3'd5};
t1 = {3'd6, 3'd6, 3'd6, 3'd2, 3'd2, 3'd2, 3'd4, 3'd4, 3'd4, 3'd6, 3'd6, 3'd6, 3'd0, 3'd0, 3'd5, 3'd5};
s0 = {1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0};
s1 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0};
//MAC result =  -10567
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd0, 3'd3, 3'd6, 3'd1, 3'd3, 3'd6, 3'd7, 3'd1, 3'd3, 3'd6, 3'd7, 3'd1, 3'd3, 3'd6, 3'd7, 3'd0};
t1 = {3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd3, 3'd3, 3'd3, 3'd3, 3'd6, 3'd6, 3'd6, 3'd6, 3'd2};
s0 = {1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1};
s1 = {1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1};
//MAC result =  -3773
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd3, 3'd4, 3'd6, 3'd0, 3'd3, 3'd4, 3'd6, 3'd0, 3'd3, 3'd4, 3'd6, 3'd0, 3'd2, 3'd4, 3'd0, 3'd2};
t1 = {3'd2, 3'd2, 3'd2, 3'd4, 3'd4, 3'd4, 3'd4, 3'd6, 3'd6, 3'd6, 3'd6, 3'd0, 3'd0, 3'd0, 3'd2, 3'd2};
s0 = {1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1};
s1 = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
//MAC result =  -7297
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd4, 3'd0, 3'd2, 3'd4, 3'd1, 3'd4, 3'd6, 3'd1, 3'd4, 3'd6, 3'd1, 3'd4, 3'd6, 3'd0, 3'd3, 3'd4};
t1 = {3'd2, 3'd6, 3'd6, 3'd6, 3'd2, 3'd2, 3'd2, 3'd4, 3'd4, 3'd4, 3'd5, 3'd5, 3'd5, 3'd0, 3'd0, 3'd0};
s0 = {1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0};
s1 = {1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1};
//MAC result =  3649
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd6, 3'd0, 3'd3, 3'd4, 3'd6, 3'd0, 3'd3, 3'd4, 3'd6, 3'd3, 3'd3, 3'd3, 3'd2, 3'd4, 3'd5, 3'd2};
t1 = {3'd0, 3'd2, 3'd2, 3'd2, 3'd2, 3'd6, 3'd6, 3'd6, 3'd6, 3'd1, 3'd5, 3'd6, 3'd0, 3'd0, 3'd0, 3'd2};
s0 = {1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
s1 = {1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
//MAC result =  -4448
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0};
t0 = {3'd4, 3'd5, 3'd2, 3'd4, 3'd5, 3'd2, 3'd4, 3'd5, 3'd0, 3'd5, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0};
t1 = {3'd2, 3'd2, 3'd4, 3'd4, 3'd4, 3'd7, 3'd7, 3'd7, 3'd0, 3'd0, 3'd5, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0};
s0 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1};
s1 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1};
//MAC result =  -4703
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd0, 3'd4, 3'd7, 3'd0, 3'd4, 3'd7, 3'd0, 3'd2, 3'd4, 3'd6, 3'd0, 3'd2, 3'd4, 3'd6, 3'd1, 3'd3};
t1 = {3'd1, 3'd1, 3'd1, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd2, 3'd6, 3'd6, 3'd6, 3'd6, 3'd2, 3'd2};
s0 = {1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0};
s1 = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0};
//MAC result =  6498
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd6, 3'd7, 3'd1, 3'd3, 3'd6, 3'd7, 3'd1, 3'd3, 3'd6, 3'd7, 3'd1, 3'd3, 3'd7, 3'd1, 3'd3, 3'd7};
t1 = {3'd2, 3'd2, 3'd4, 3'd4, 3'd4, 3'd4, 3'd5, 3'd5, 3'd5, 3'd5, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1};
s0 = {1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1};
s1 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
//MAC result =  -3202
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd1, 3'd3, 3'd7, 3'd0, 3'd2, 3'd4, 3'd0, 3'd2, 3'd4, 3'd0, 3'd2, 3'd4, 3'd0, 3'd2, 3'd4, 3'd0};
t1 = {3'd3, 3'd3, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd4, 3'd4, 3'd4, 3'd7, 3'd7, 3'd7, 3'd2};
s0 = {1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1};
s1 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0};
//MAC result =  469
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd2, 3'd0, 3'd2, 3'd0, 3'd2, 3'd1, 3'd7, 3'd1, 3'd7, 3'd1, 3'd7, 3'd0, 3'd2, 3'd0, 3'd2, 3'd0};
t1 = {3'd2, 3'd4, 3'd4, 3'd6, 3'd6, 3'd0, 3'd0, 3'd5, 3'd5, 3'd7, 3'd7, 3'd1, 3'd1, 3'd4, 3'd4, 3'd6};
s0 = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0};
s1 = {1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1};
//MAC result =  12312
//-------------------------------
#5;

in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
t0 = {3'd2, 3'd0, 3'd5, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0};
t1 = {3'd6, 3'd0, 3'd0, 3'd5, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0};
s0 = {1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
s1 = {1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
//MAC result =  1217
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd1, 3'd6, 3'd1, 3'd6, 3'd1, 3'd6, 3'd0, 3'd2, 3'd0, 3'd2, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2};
t1 = {3'd0, 3'd0, 3'd5, 3'd5, 3'd6, 3'd6, 3'd1, 3'd1, 3'd4, 3'd4, 3'd0, 3'd3, 3'd5, 3'd6, 3'd2, 3'd2};
s0 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1};
s1 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0};
//MAC result =  6295
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd6, 3'd0, 3'd2, 3'd6, 3'd4, 3'd4, 3'd4, 3'd4, 3'd0, 3'd1, 3'd6, 3'd0, 3'd1, 3'd6, 3'd0, 3'd1};
t1 = {3'd2, 3'd4, 3'd4, 3'd4, 3'd1, 3'd3, 3'd4, 3'd7, 3'd0, 3'd0, 3'd0, 3'd2, 3'd2, 3'd2, 3'd7, 3'd7};
s0 = {1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
s1 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1};
//MAC result =  -3265
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd6, 3'd0, 3'd3, 3'd4, 3'd6, 3'd0, 3'd3, 3'd4, 3'd6, 3'd0, 3'd3, 3'd6, 3'd0, 3'd3, 3'd6, 3'd0};
t1 = {3'd7, 3'd0, 3'd0, 3'd0, 3'd0, 3'd4, 3'd4, 3'd4, 3'd4, 3'd5, 3'd5, 3'd5, 3'd6, 3'd6, 3'd6, 3'd0};
s0 = {1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1};
s1 = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1};
//MAC result =  -12966
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
t0 = {3'd5, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0};
t1 = {3'd0, 3'd5, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0};
s0 = {1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
s1 = {1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
//MAC result =  992
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd1, 3'd3, 3'd5, 3'd7, 3'd1, 3'd3, 3'd5, 3'd7, 3'd1, 3'd3, 3'd5, 3'd7, 3'd0, 3'd2, 3'd4, 3'd0};
t1 = {3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd2, 3'd2, 3'd2, 3'd5, 3'd5, 3'd5, 3'd5, 3'd0, 3'd0, 3'd0, 3'd4};
s0 = {1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
s1 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
//MAC result =  -2515
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd2, 3'd4, 3'd0, 3'd2, 3'd4, 3'd1, 3'd6, 3'd1, 3'd6, 3'd1, 3'd6, 3'd6, 3'd6, 3'd1, 3'd5, 3'd7};
t1 = {3'd4, 3'd4, 3'd6, 3'd6, 3'd6, 3'd3, 3'd3, 3'd5, 3'd5, 3'd6, 3'd6, 3'd4, 3'd6, 3'd3, 3'd3, 3'd3};
s0 = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1};
s1 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0};
//MAC result =  -1920
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd1, 3'd5, 3'd7, 3'd1, 3'd5, 3'd7, 3'd2, 3'd4, 3'd6, 3'd2, 3'd4, 3'd6, 3'd2, 3'd4, 3'd6, 3'd0};
t1 = {3'd4, 3'd4, 3'd4, 3'd6, 3'd6, 3'd6, 3'd1, 3'd1, 3'd1, 3'd4, 3'd4, 3'd4, 3'd5, 3'd5, 3'd5, 3'd0};
s0 = {1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
s1 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
//MAC result =  -3319
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd3, 3'd5, 3'd7, 3'd0, 3'd3, 3'd5, 3'd7, 3'd0, 3'd3, 3'd5, 3'd7, 3'd0, 3'd3, 3'd4, 3'd6, 3'd0};
t1 = {3'd0, 3'd0, 3'd0, 3'd3, 3'd3, 3'd3, 3'd3, 3'd6, 3'd6, 3'd6, 3'd6, 3'd1, 3'd1, 3'd1, 3'd1, 3'd6};
s0 = {1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1};
s1 = {1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
//MAC result =  5966
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
t0 = {3'd3, 3'd4, 3'd6, 3'd0, 3'd3, 3'd4, 3'd6, 3'd0, 3'd5, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0};
t1 = {3'd6, 3'd6, 3'd6, 3'd7, 3'd7, 3'd7, 3'd7, 3'd0, 3'd0, 3'd5, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0};
s0 = {1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
s1 = {1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
//MAC result =  5697
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd4, 3'd4, 3'd4, 3'd2, 3'd5, 3'd2, 3'd5, 3'd2, 3'd5, 3'd2, 3'd4, 3'd6, 3'd2, 3'd4, 3'd6, 3'd2};
t1 = {3'd1, 3'd5, 3'd6, 3'd0, 3'd0, 3'd2, 3'd2, 3'd7, 3'd7, 3'd0, 3'd0, 3'd0, 3'd2, 3'd2, 3'd2, 3'd3};
s0 = {1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
s1 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
//MAC result =  4616
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd4, 3'd6, 3'd2, 3'd4, 3'd6, 3'd2, 3'd4, 3'd6, 3'd2, 3'd4, 3'd6, 3'd1, 3'd2, 3'd4, 3'd1, 3'd2};
t1 = {3'd3, 3'd3, 3'd7, 3'd7, 3'd7, 3'd1, 3'd1, 3'd1, 3'd7, 3'd7, 3'd7, 3'd0, 3'd0, 3'd0, 3'd2, 3'd2};
s0 = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
s1 = {1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1};
//MAC result =  20698
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd4, 3'd1, 3'd2, 3'd4, 3'd1, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd5, 3'd0, 3'd2, 3'd3, 3'd5, 3'd0};
t1 = {3'd2, 3'd5, 3'd5, 3'd5, 3'd6, 3'd6, 3'd6, 3'd4, 3'd4, 3'd7, 3'd7, 3'd0, 3'd0, 3'd0, 3'd0, 3'd2};
s0 = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
s1 = {1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
//MAC result =  -5471
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd2, 3'd3, 3'd5, 3'd0, 3'd2, 3'd3, 3'd5, 3'd0, 3'd2, 3'd6, 3'd0, 3'd2, 3'd6, 3'd0, 3'd2, 3'd6};
t1 = {3'd2, 3'd2, 3'd2, 3'd5, 3'd5, 3'd5, 3'd5, 3'd0, 3'd0, 3'd0, 3'd2, 3'd2, 3'd2, 3'd6, 3'd6, 3'd6};
s0 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0};
s1 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0};
//MAC result =  5097
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
t0 = {3'd0, 3'd5, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0};
t1 = {3'd0, 3'd0, 3'd5, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0};
s0 = {1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
s1 = {1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
//MAC result =  993
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd1, 3'd2, 3'd6, 3'd1, 3'd2, 3'd6, 3'd1, 3'd2, 3'd6, 3'd1, 3'd2, 3'd6, 3'd1, 3'd4, 3'd7, 3'd1};
t1 = {3'd0, 3'd0, 3'd0, 3'd3, 3'd3, 3'd3, 3'd5, 3'd5, 3'd5, 3'd6, 3'd6, 3'd6, 3'd0, 3'd0, 3'd0, 3'd4};
s0 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0};
s1 = {1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0};
//MAC result =  -6088
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd4, 3'd7, 3'd0, 3'd4, 3'd0, 3'd4, 3'd0, 3'd1, 3'd5, 3'd7, 3'd0, 3'd1, 3'd5, 3'd7, 3'd0, 3'd1};
t1 = {3'd4, 3'd4, 3'd0, 3'd0, 3'd3, 3'd3, 3'd1, 3'd1, 3'd1, 3'd1, 3'd5, 3'd5, 3'd5, 3'd5, 3'd7, 3'd7};
s0 = {1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0};
s1 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1};
//MAC result =  -5101
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd5, 3'd7, 3'd0, 3'd2, 3'd5, 3'd0, 3'd2, 3'd5, 3'd0, 3'd2, 3'd5, 3'd1, 3'd3, 3'd6, 3'd7, 3'd1};
t1 = {3'd7, 3'd7, 3'd1, 3'd1, 3'd1, 3'd4, 3'd4, 3'd4, 3'd6, 3'd6, 3'd6, 3'd1, 3'd1, 3'd1, 3'd1, 3'd3};
s0 = {1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0};
s1 = {1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
//MAC result =  14574
//-------------------------------
#5;

in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd3, 3'd6, 3'd7, 3'd1, 3'd3, 3'd6, 3'd7, 3'd0, 3'd2, 3'd0, 3'd2, 3'd0, 3'd2, 3'd0, 3'd2, 3'd6};
t1 = {3'd3, 3'd3, 3'd3, 3'd6, 3'd6, 3'd6, 3'd6, 3'd2, 3'd2, 3'd5, 3'd5, 3'd6, 3'd6, 3'd1, 3'd1, 3'd1};
s0 = {1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1};
s1 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
//MAC result =  -4302
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
t0 = {3'd0, 3'd2, 3'd6, 3'd0, 3'd5, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0};
t1 = {3'd6, 3'd6, 3'd6, 3'd0, 3'd0, 3'd5, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0};
s0 = {1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
s1 = {1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
//MAC result =  -2943
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd0, 3'd2, 3'd4, 3'd6, 3'd0, 3'd2, 3'd4, 3'd6, 3'd0, 3'd2, 3'd4, 3'd6, 3'd0, 3'd3, 3'd4, 3'd7};
t1 = {3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd2, 3'd2, 3'd2, 3'd6, 3'd6, 3'd6, 3'd6, 3'd0, 3'd0, 3'd0, 3'd0};
s0 = {1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1};
s1 = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
//MAC result =  -4648
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd0, 3'd3, 3'd4, 3'd7, 3'd0, 3'd3, 3'd4, 3'd7, 3'd0, 3'd3, 3'd4, 3'd7, 3'd3, 3'd7, 3'd3, 3'd7};
t1 = {3'd3, 3'd3, 3'd3, 3'd3, 3'd4, 3'd4, 3'd4, 3'd4, 3'd6, 3'd6, 3'd6, 3'd6, 3'd3, 3'd3, 3'd5, 3'd5};
s0 = {1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1};
s1 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0};
//MAC result =  -12120
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd3, 3'd7, 3'd0, 3'd5, 3'd6, 3'd0, 3'd5, 3'd6, 3'd0, 3'd5, 3'd6, 3'd0, 3'd3, 3'd6, 3'd0, 3'd3};
t1 = {3'd6, 3'd6, 3'd2, 3'd2, 3'd2, 3'd5, 3'd5, 3'd5, 3'd7, 3'd7, 3'd7, 3'd0, 3'd0, 3'd0, 3'd2, 3'd2};
s0 = {1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1};
s1 = {1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
//MAC result =  -1159
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd6, 3'd0, 3'd3, 3'd6, 3'd0, 3'd3, 3'd6, 3'd3, 3'd7, 3'd3, 3'd7, 3'd3, 3'd7, 3'd0, 3'd2, 3'd5};
t1 = {3'd2, 3'd4, 3'd4, 3'd4, 3'd7, 3'd7, 3'd7, 3'd0, 3'd0, 3'd4, 3'd4, 3'd6, 3'd6, 3'd0, 3'd0, 3'd0};
s0 = {1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0};
s1 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
//MAC result =  -1997
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd6, 3'd0, 3'd2, 3'd5, 3'd6, 3'd0, 3'd2, 3'd5, 3'd6, 3'd0, 3'd2, 3'd5, 3'd6, 3'd2, 3'd6, 3'd2};
t1 = {3'd0, 3'd2, 3'd2, 3'd2, 3'd2, 3'd3, 3'd3, 3'd3, 3'd3, 3'd5, 3'd5, 3'd5, 3'd5, 3'd0, 3'd0, 3'd2};
s0 = {1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1};
s1 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0};
//MAC result =  4120
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
t0 = {3'd6, 3'd2, 3'd6, 3'd0, 3'd5, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0};
t1 = {3'd2, 3'd4, 3'd4, 3'd0, 3'd0, 3'd5, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0};
s0 = {1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
s1 = {1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
//MAC result =  1793
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd1, 3'd4, 3'd1, 3'd4, 3'd0, 3'd2, 3'd4, 3'd6, 3'd0, 3'd2, 3'd4, 3'd6, 3'd2, 3'd5, 3'd6, 3'd2};
t1 = {3'd4, 3'd4, 3'd7, 3'd7, 3'd4, 3'd4, 3'd4, 3'd4, 3'd7, 3'd7, 3'd7, 3'd7, 3'd0, 3'd0, 3'd0, 3'd4};
s0 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0};
s1 = {1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
//MAC result =  -11212
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd5, 3'd6, 3'd2, 3'd5, 3'd6, 3'd0, 3'd2, 3'd7, 3'd0, 3'd2, 3'd7, 3'd0, 3'd2, 3'd7, 3'd0, 3'd2};
t1 = {3'd4, 3'd4, 3'd5, 3'd5, 3'd5, 3'd0, 3'd0, 3'd0, 3'd2, 3'd2, 3'd2, 3'd4, 3'd4, 3'd4, 3'd6, 3'd6};
s0 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1};
s1 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1};
//MAC result =  6553
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd7, 3'd0, 3'd1, 3'd3, 3'd5, 3'd0, 3'd1, 3'd3, 3'd5, 3'd0, 3'd3, 3'd4, 3'd6, 3'd0, 3'd3, 3'd4};
t1 = {3'd6, 3'd1, 3'd1, 3'd1, 3'd1, 3'd6, 3'd6, 3'd6, 3'd6, 3'd0, 3'd0, 3'd0, 3'd0, 3'd5, 3'd5, 3'd5};
s0 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0};
s1 = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1};
//MAC result =  -11679
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0};
t0 = {3'd6, 3'd1, 3'd2, 3'd1, 3'd2, 3'd3, 3'd4, 3'd6, 3'd3, 3'd4, 3'd6, 3'd0, 3'd5, 3'd0, 3'd5, 3'd0};
t1 = {3'd5, 3'd0, 3'd0, 3'd6, 3'd6, 3'd3, 3'd3, 3'd3, 3'd4, 3'd4, 3'd4, 3'd0, 3'd0, 3'd5, 3'd5, 3'd0};
s0 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1};
s1 = {1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1};
//MAC result =  -2821
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd0, 3'd1, 3'd2, 3'd5, 3'd0, 3'd1, 3'd2, 3'd5, 3'd0, 3'd1, 3'd2, 3'd5, 3'd0, 3'd1, 3'd2, 3'd5};
t1 = {3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd2, 3'd2, 3'd2, 3'd4, 3'd4, 3'd4, 3'd4, 3'd6, 3'd6, 3'd6, 3'd6};
s0 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
s1 = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1};
//MAC result =  -2067
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd0, 3'd3, 3'd6, 3'd0, 3'd3, 3'd6, 3'd0, 3'd3, 3'd6, 3'd2, 3'd7, 3'd2, 3'd7, 3'd1, 3'd3, 3'd5};
t1 = {3'd0, 3'd0, 3'd0, 3'd2, 3'd2, 3'd2, 3'd4, 3'd4, 3'd4, 3'd2, 3'd2, 3'd3, 3'd3, 3'd0, 3'd0, 3'd0};
s0 = {1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0};
s1 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
//MAC result =  -2073
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd6, 3'd1, 3'd3, 3'd5, 3'd6, 3'd1, 3'd3, 3'd5, 3'd6, 3'd1, 3'd3, 3'd5, 3'd6, 3'd1, 3'd4, 3'd1};
t1 = {3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd3, 3'd3, 3'd3, 3'd3, 3'd6, 3'd6, 3'd6, 3'd6, 3'd2, 3'd2, 3'd6};
s0 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1};
s1 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1};
//MAC result =  8092
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd4, 3'd1, 3'd2, 3'd4, 3'd1, 3'd2, 3'd4, 3'd1, 3'd2, 3'd4, 3'd0, 3'd3, 3'd0, 3'd3, 3'd0, 3'd3};
t1 = {3'd6, 3'd1, 3'd1, 3'd1, 3'd2, 3'd2, 3'd2, 3'd6, 3'd6, 3'd6, 3'd0, 3'd0, 3'd5, 3'd5, 3'd7, 3'd7};
s0 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0};
s1 = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1};
//MAC result =  -3243
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0};
t0 = {3'd0, 3'd2, 3'd4, 3'd0, 3'd2, 3'd4, 3'd0, 3'd2, 3'd4, 3'd0, 3'd5, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0};
t1 = {3'd1, 3'd1, 3'd1, 3'd2, 3'd2, 3'd2, 3'd5, 3'd5, 3'd5, 3'd0, 3'd0, 3'd5, 3'd5, 3'd0, 3'd0, 3'd0};
s0 = {1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1};
s1 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1};
//MAC result =  467
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd3, 3'd3, 3'd0, 3'd2, 3'd6, 3'd0, 3'd2, 3'd6, 3'd0, 3'd2, 3'd6, 3'd2, 3'd4, 3'd6, 3'd2, 3'd4};
t1 = {3'd4, 3'd7, 3'd0, 3'd0, 3'd0, 3'd2, 3'd2, 3'd2, 3'd7, 3'd7, 3'd7, 3'd1, 3'd1, 3'd1, 3'd5, 3'd5};
s0 = {1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0};
s1 = {1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
//MAC result =  -8719
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};

t0 = {3'd6, 3'd2, 3'd4, 3'd6, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd1, 3'd0, 3'd3, 3'd6, 3'd2, 3'd4, 3'd2};
t1 = {3'd5, 3'd6, 3'd6, 3'd6, 3'd0, 3'd0, 3'd2, 3'd2, 3'd6, 3'd6, 3'd6, 3'd6, 3'd6, 3'd1, 3'd1, 3'd3};
s0 = {1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0};
s1 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0};
//MAC result =  -8313
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd4, 3'd2, 3'd4, 3'd2, 3'd4, 3'd0, 3'd2, 3'd5, 3'd0, 3'd2, 3'd5, 3'd0, 3'd2, 3'd5, 3'd3, 3'd6};
t1 = {3'd3, 3'd4, 3'd4, 3'd7, 3'd7, 3'd2, 3'd2, 3'd2, 3'd5, 3'd5, 3'd5, 3'd6, 3'd6, 3'd6, 3'd1, 3'd1};
s0 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
s1 = {1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1};
//MAC result =  5924
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
t0 = {3'd3, 3'd6, 3'd0, 3'd5, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0};
t1 = {3'd6, 3'd6, 3'd0, 3'd0, 3'd5, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0};
s0 = {1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
s1 = {1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
//MAC result =  5601
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd0, 3'd2, 3'd4, 3'd6, 3'd0, 3'd2, 3'd4, 3'd6, 3'd0, 3'd2, 3'd4, 3'd6, 3'd0, 3'd2, 3'd4, 3'd6};
t1 = {3'd0, 3'd0, 3'd0, 3'd0, 3'd3, 3'd3, 3'd3, 3'd3, 3'd5, 3'd5, 3'd5, 3'd5, 3'd6, 3'd6, 3'd6, 3'd6};
s0 = {1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1};
s1 = {1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
//MAC result =  6675
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd3, 3'd5, 3'd6, 3'd3, 3'd5, 3'd6, 3'd3, 3'd5, 3'd6, 3'd3, 3'd5, 3'd6, 3'd0, 3'd1, 3'd5, 3'd2};
t1 = {3'd1, 3'd1, 3'd1, 3'd2, 3'd2, 3'd2, 3'd4, 3'd4, 3'd4, 3'd5, 3'd5, 3'd5, 3'd4, 3'd4, 3'd4, 3'd1};
s0 = {1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0};
s1 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1};
//MAC result =  -1608
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd3, 3'd7, 3'd2, 3'd3, 3'd7, 3'd2, 3'd3, 3'd7, 3'd2, 3'd5, 3'd2, 3'd5, 3'd2, 3'd5, 3'd2, 3'd3};
t1 = {3'd1, 3'd1, 3'd4, 3'd4, 3'd4, 3'd6, 3'd6, 3'd6, 3'd0, 3'd0, 3'd4, 3'd4, 3'd5, 3'd5, 3'd2, 3'd2};
s0 = {1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
s1 = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
//MAC result =  -3516
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd6, 3'd2, 3'd3, 3'd6, 3'd2, 3'd3, 3'd6, 3'd0, 3'd3, 3'd4, 3'd6, 3'd0, 3'd3, 3'd4, 3'd6, 3'd0};
t1 = {3'd2, 3'd5, 3'd5, 3'd5, 3'd6, 3'd6, 3'd6, 3'd1, 3'd1, 3'd1, 3'd1, 3'd2, 3'd2, 3'd2, 3'd2, 3'd4};
s0 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
s1 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1};
//MAC result =  7458
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0};
t0 = {3'd3, 3'd4, 3'd6, 3'd1, 3'd6, 3'd1, 3'd6, 3'd1, 3'd6, 3'd0, 3'd5, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0};
t1 = {3'd4, 3'd4, 3'd4, 3'd0, 3'd0, 3'd3, 3'd3, 3'd7, 3'd7, 3'd0, 3'd0, 3'd5, 3'd5, 3'd0, 3'd0, 3'd0};
s0 = {1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1};
s1 = {1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1};
//MAC result =  -7825
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd1, 3'd4, 3'd7, 3'd1, 3'd4, 3'd7, 3'd1, 3'd4, 3'd7, 3'd2, 3'd2, 3'd2, 3'd1, 3'd4, 3'd6, 3'd1};
t1 = {3'd1, 3'd1, 3'd1, 3'd4, 3'd4, 3'd4, 3'd7, 3'd7, 3'd7, 3'd0, 3'd2, 3'd5, 3'd3, 3'd3, 3'd3, 3'd5};
s0 = {1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1};
s1 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
//MAC result =  12992
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd4, 3'd6, 3'd1, 3'd4, 3'd6, 3'd0, 3'd2, 3'd5, 3'd0, 3'd2, 3'd5, 3'd0, 3'd3, 3'd4, 3'd7, 3'd0};
t1 = {3'd5, 3'd5, 3'd6, 3'd6, 3'd6, 3'd4, 3'd4, 3'd4, 3'd7, 3'd7, 3'd7, 3'd0, 3'd0, 3'd0, 3'd0, 3'd3};
s0 = {1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1};
s1 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1};
//MAC result =  10703
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd3, 3'd4, 3'd7, 3'd0, 3'd3, 3'd4, 3'd7, 3'd0, 3'd7, 3'd0, 3'd7, 3'd0, 3'd7, 3'd2, 3'd2, 3'd2};
t1 = {3'd3, 3'd3, 3'd3, 3'd7, 3'd7, 3'd7, 3'd7, 3'd2, 3'd2, 3'd3, 3'd3, 3'd5, 3'd5, 3'd0, 3'd3, 3'd4};
s0 = {1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0};
s1 = {1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1};
//MAC result =  -7112
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd0, 3'd3, 3'd5, 3'd6, 3'd0, 3'd3, 3'd5, 3'd6, 3'd0, 3'd3, 3'd5, 3'd6, 3'd0, 3'd3, 3'd5, 3'd6};
t1 = {3'd0, 3'd0, 3'd0, 3'd0, 3'd3, 3'd3, 3'd3, 3'd3, 3'd5, 3'd5, 3'd5, 3'd5, 3'd6, 3'd6, 3'd6, 3'd6};
s0 = {1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1};
s1 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
//MAC result =  -4095
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
t0 = {3'd0, 3'd5, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0};
t1 = {3'd0, 3'd0, 3'd5, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0};
s0 = {1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
s1 = {1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
//MAC result =  993
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd3, 3'd5, 3'd6, 3'd3, 3'd5, 3'd6, 3'd3, 3'd5, 3'd6, 3'd0, 3'd4, 3'd7, 3'd0, 3'd4, 3'd7, 3'd0};
t1 = {3'd0, 3'd0, 3'd0, 3'd5, 3'd5, 3'd5, 3'd6, 3'd6, 3'd6, 3'd2, 3'd2, 3'd2, 3'd4, 3'd4, 3'd4, 3'd6};
s0 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0};
s1 = {1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1};
//MAC result =  11148
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd4, 3'd7, 3'd0, 3'd4, 3'd7, 3'd0, 3'd4, 3'd7, 3'd1, 3'd1, 3'd3, 3'd5, 3'd6, 3'd1, 3'd3, 3'd5};
t1 = {3'd6, 3'd6, 3'd0, 3'd0, 3'd0, 3'd4, 3'd4, 3'd4, 3'd7, 3'd2, 3'd2, 3'd2, 3'd2, 3'd5, 3'd5, 3'd5};
s0 = {1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
s1 = {1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1};
//MAC result =  8169
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd6, 3'd0, 3'd3, 3'd6, 3'd0, 3'd3, 3'd6, 3'd0, 3'd3, 3'd6, 3'd0, 3'd1, 3'd7, 3'd0, 3'd1, 3'd7};
t1 = {3'd5, 3'd0, 3'd0, 3'd0, 3'd4, 3'd4, 3'd4, 3'd7, 3'd7, 3'd7, 3'd0, 3'd0, 3'd0, 3'd3, 3'd3, 3'd3};
s0 = {1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1};
s1 = {1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0};
//MAC result =  3518
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0};
t0 = {3'd0, 3'd1, 3'd7, 3'd0, 3'd3, 3'd5, 3'd0, 3'd3, 3'd5, 3'd0, 3'd5, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0};
t1 = {3'd4, 3'd4, 3'd4, 3'd1, 3'd1, 3'd1, 3'd4, 3'd4, 3'd4, 3'd0, 3'd0, 3'd5, 3'd5, 3'd0, 3'd0, 3'd0};
s0 = {1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1};
s1 = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1};
//MAC result =  3535
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd0, 3'd2, 3'd7, 3'd0, 3'd2, 3'd7, 3'd0, 3'd2, 3'd7, 3'd5, 3'd5, 3'd4, 3'd7, 3'd4, 3'd7, 3'd4};
t1 = {3'd1, 3'd1, 3'd1, 3'd3, 3'd3, 3'd3, 3'd4, 3'd4, 3'd4, 3'd3, 3'd5, 3'd1, 3'd1, 3'd4, 3'd4, 3'd7};
s0 = {1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1};
s1 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0};
//MAC result =  -6494
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd7, 3'd0, 3'd5, 3'd0, 3'd5, 3'd0, 3'd5, 3'd0, 3'd5, 3'd0, 3'd7, 3'd0, 3'd7, 3'd0, 3'd7, 3'd0};
t1 = {3'd7, 3'd1, 3'd1, 3'd2, 3'd2, 3'd4, 3'd4, 3'd5, 3'd5, 3'd1, 3'd1, 3'd4, 3'd4, 3'd7, 3'd7, 3'd1};
s0 = {1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1};
s1 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0};
//MAC result =  4086
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd3, 3'd4, 3'd0, 3'd3, 3'd4, 3'd0, 3'd3, 3'd4, 3'd0, 3'd3, 3'd6, 3'd0, 3'd3, 3'd6, 3'd0, 3'd3};
t1 = {3'd1, 3'd1, 3'd5, 3'd5, 3'd5, 3'd7, 3'd7, 3'd7, 3'd0, 3'd0, 3'd0, 3'd2, 3'd2, 3'd2, 3'd4, 3'd4};
s0 = {1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0};
s1 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
//MAC result =  939
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0};

t0 = {3'd6, 3'd1, 3'd4, 3'd5, 3'd6, 3'd1, 3'd4, 3'd5, 3'd6, 3'd0, 3'd5, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0};
t1 = {3'd4, 3'd4, 3'd4, 3'd4, 3'd4, 3'd5, 3'd5, 3'd5, 3'd5, 3'd0, 3'd0, 3'd5, 3'd5, 3'd0, 3'd0, 3'd0};
s0 = {1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1};
s1 = {1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1};
//MAC result =  7457
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd1, 3'd1, 3'd1, 3'd1, 3'd0, 3'd2, 3'd4, 3'd0, 3'd2, 3'd4, 3'd0, 3'd2, 3'd4, 3'd0, 3'd2, 3'd4};
t1 = {3'd1, 3'd2, 3'd4, 3'd6, 3'd0, 3'd0, 3'd0, 3'd2, 3'd2, 3'd2, 3'd5, 3'd5, 3'd5, 3'd7, 3'd7, 3'd7};
s0 = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1};
s1 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1};
//MAC result =  1011
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
t0 = {3'd0, 3'd6, 3'd0, 3'd6, 3'd2, 3'd3, 3'd5, 3'd2, 3'd3, 3'd5, 3'd2, 3'd3, 3'd5, 3'd2, 3'd4, 3'd7};
t1 = {3'd1, 3'd1, 3'd5, 3'd5, 3'd0, 3'd0, 3'd0, 3'd4, 3'd4, 3'd4, 3'd7, 3'd7, 3'd7, 3'd2, 3'd2, 3'd2};
s0 = {1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0};
s1 = {1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
//MAC result =  3486
//-------------------------------
#5;
in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0};
t0 = {3'd2, 3'd4, 3'd7, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd5, 3'd0, 3'd5, 3'd0, 3'd0};
t1 = {3'd5, 3'd5, 3'd5, 3'd0, 3'd4, 3'd6, 3'd1, 3'd3, 3'd4, 3'd6, 3'd0, 3'd0, 3'd5, 3'd5, 3'd0, 3'd0};
s0 = {1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1};
s1 = {1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1};
//MAC result =  -2598


    end
    
endmodule
