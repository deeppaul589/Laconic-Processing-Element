`timescale 1ns / 1ps

module tb();
    
    reg [15:0] in_applied;
    reg [47:0] t0;
    reg [47:0] t1;
    reg [15:0] s0;
    reg [15:0] s1;
    
    wire signed [21:0] result;
    
    core uut(
    
        .in_applied(in_applied),
        .t0(t0),
        .t1(t1),
        .s0(s0),
        .s1(s1),
        .out_value(result)
    
    );
    
    
    
    initial begin
        
        #5; 
        //210
        in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0};
        
        t0 = {3'd5, 3'd5, 3'd5, 3'd3, 3'd3, 3'd3, 3'd2, 3'd2, 3'd2, 3'd1, 3'd1, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0};
        // A = (2^5-2^3+2^2+2^1)
        t1 = {3'd2, 3'd1, 3'd0, 3'd2, 3'd1, 3'd0, 3'd2, 3'd1, 3'd0, 3'd2, 3'd1, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0};
        // B = (2^2+2^1+2^0)
        
        s0 = {1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
        s1 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
        
		//-------------------------------
		#5;
		in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
		t0 = {3'd0, 3'd1, 3'd4, 3'd0, 3'd1, 3'd4, 3'd0, 3'd1, 3'd4, 3'd0, 3'd0, 3'd0, 3'd7, 3'd0, 3'd4, 3'd7};
		t1 = {3'd0, 3'd0, 3'd0, 3'd2, 3'd2, 3'd2, 3'd4, 3'd4, 3'd4, 3'd1, 3'd2, 3'd6, 3'd3, 3'd0, 3'd0, 3'd0};
		s0 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0};
		s1 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0};
		//MAC result =  856
		//-------------------------------
		#5;
		in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
		t0 = {3'd0, 3'd4, 3'd7, 3'd0, 3'd4, 3'd7, 3'd1, 3'd4, 3'd1, 3'd4, 3'd1, 3'd4, 3'd7, 3'd7, 3'd7, 3'd2};
		t1 = {3'd1, 3'd1, 3'd1, 3'd4, 3'd4, 3'd4, 3'd0, 3'd0, 3'd2, 3'd2, 3'd5, 3'd5, 3'd0, 3'd4, 3'd6, 3'd0};
		s0 = {1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0};
		s1 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1};
		//MAC result =  8752
		//-------------------------------
		#5;
		in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
		t0 = {3'd3, 3'd2, 3'd3, 3'd7, 3'd7, 3'd7, 3'd7, 3'd7, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0};
		t1 = {3'd0, 3'd5, 3'd5, 3'd0, 3'd3, 3'd4, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0};
		s0 = {1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
		s1 = {1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
		//MAC result =  -6792
		//-------------------------------
		#5;
		in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
		t0 = {3'd0, 3'd1, 3'd4, 3'd0, 3'd1, 3'd4, 3'd0, 3'd1, 3'd4, 3'd0, 3'd0, 3'd0, 3'd7, 3'd0, 3'd4, 3'd7};
		t1 = {3'd0, 3'd0, 3'd0, 3'd2, 3'd2, 3'd2, 3'd4, 3'd4, 3'd4, 3'd1, 3'd2, 3'd6, 3'd3, 3'd0, 3'd0, 3'd0};
		s0 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0};
		s1 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0};
		//MAC result =  856
		//-------------------------------
		#5;
		in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
		t0 = {3'd0, 3'd4, 3'd7, 3'd0, 3'd4, 3'd7, 3'd1, 3'd4, 3'd1, 3'd4, 3'd1, 3'd4, 3'd7, 3'd7, 3'd7, 3'd2};
		t1 = {3'd1, 3'd1, 3'd1, 3'd4, 3'd4, 3'd4, 3'd0, 3'd0, 3'd2, 3'd2, 3'd5, 3'd5, 3'd0, 3'd4, 3'd6, 3'd0};
		s0 = {1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0};
		s1 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1};
		//MAC result =  8752
		//-------------------------------
		#5;
		in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
		t0 = {3'd3, 3'd2, 3'd3, 3'd7, 3'd7, 3'd7, 3'd0, 3'd5, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0};
		t1 = {3'd0, 3'd5, 3'd5, 3'd0, 3'd3, 3'd4, 3'd0, 3'd0, 3'd5, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0};
		s0 = {1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
		s1 = {1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
		//MAC result =  -1607
		//-------------------------------
		#5;
		in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
		t0 = {3'd0, 3'd1, 3'd4, 3'd0, 3'd1, 3'd4, 3'd0, 3'd1, 3'd4, 3'd0, 3'd0, 3'd0, 3'd7, 3'd0, 3'd4, 3'd7};
		t1 = {3'd0, 3'd0, 3'd0, 3'd2, 3'd2, 3'd2, 3'd4, 3'd4, 3'd4, 3'd1, 3'd2, 3'd6, 3'd3, 3'd0, 3'd0, 3'd0};
		s0 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0};
		s1 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0};
		//MAC result =  -1192
		//-------------------------------
		#5;
		in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
		t0 = {3'd0, 3'd4, 3'd7, 3'd0, 3'd4, 3'd7, 3'd1, 3'd4, 3'd1, 3'd4, 3'd1, 3'd4, 3'd7, 3'd7, 3'd7, 3'd2};
		t1 = {3'd1, 3'd1, 3'd1, 3'd4, 3'd4, 3'd4, 3'd0, 3'd0, 3'd2, 3'd2, 3'd5, 3'd5, 3'd0, 3'd4, 3'd6, 3'd0};
		s0 = {1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0};
		s1 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1};
		//MAC result =  8752
		//-------------------------------
		#5;
		in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
		t0 = {3'd3, 3'd2, 3'd3, 3'd7, 3'd7, 3'd7, 3'd0, 3'd5, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0};
		t1 = {3'd0, 3'd5, 3'd5, 3'd0, 3'd3, 3'd4, 3'd0, 3'd0, 3'd5, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0};
		s0 = {1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
		s1 = {1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
		//MAC result =  -1607
		//-------------------------------
		#5;
		in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
		t0 = {3'd0, 3'd3, 3'd4, 3'd7, 3'd0, 3'd3, 3'd4, 3'd7, 3'd0, 3'd3, 3'd4, 3'd7, 3'd1, 3'd3, 3'd1, 3'd3};
		t1 = {3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd2, 3'd2, 3'd2, 3'd4, 3'd4, 3'd4, 3'd4, 3'd0, 3'd0, 3'd3, 3'd3};
		s0 = {1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
		s1 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1};
		//MAC result =  -1379
		//-------------------------------
		#5;
		in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
		t0 = {3'd1, 3'd3, 3'd2, 3'd4, 3'd0, 3'd1, 3'd3, 3'd0, 3'd1, 3'd3, 3'd0, 3'd1, 3'd3, 3'd1, 3'd4, 3'd1};
		t1 = {3'd6, 3'd6, 3'd3, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd4, 3'd4, 3'd4, 3'd0, 3'd0, 3'd2};
		s0 = {1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
		s1 = {1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1};
		//MAC result =  -553
		//-------------------------------
		#5;
		in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
		t0 = {3'd4, 3'd1, 3'd4, 3'd7, 3'd7, 3'd7, 3'd2, 3'd3, 3'd2, 3'd3, 3'd7, 3'd7, 3'd7, 3'd0, 3'd5, 3'd0};
		t1 = {3'd2, 3'd5, 3'd5, 3'd0, 3'd4, 3'd6, 3'd0, 3'd0, 3'd5, 3'd5, 3'd0, 3'd3, 3'd4, 3'd0, 3'd0, 3'd5};
		s0 = {1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1};
		s1 = {1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0};
		//MAC result =  4149
		//-------------------------------
		#5;
		in_applied = {1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
		t0 = {3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0};
		t1 = {3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0};
		s0 = {1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
		s1 = {1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
		//MAC result =  1024
		//-------------------------------
		#5;
		in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
		t0 = {3'd0, 3'd3, 3'd4, 3'd7, 3'd0, 3'd3, 3'd4, 3'd7, 3'd0, 3'd3, 3'd4, 3'd7, 3'd1, 3'd3, 3'd1, 3'd3};
		t1 = {3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd2, 3'd2, 3'd2, 3'd4, 3'd4, 3'd4, 3'd4, 3'd0, 3'd0, 3'd3, 3'd3};
		s0 = {1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
		s1 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1};
		//MAC result =  -1379
		//-------------------------------
		#5;
		in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
		t0 = {3'd1, 3'd3, 3'd2, 3'd4, 3'd0, 3'd1, 3'd3, 3'd0, 3'd1, 3'd3, 3'd0, 3'd1, 3'd3, 3'd1, 3'd4, 3'd1};
		t1 = {3'd6, 3'd6, 3'd3, 3'd3, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd4, 3'd4, 3'd4, 3'd0, 3'd0, 3'd2};
		s0 = {1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
		s1 = {1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1};
		//MAC result =  -553
		//-------------------------------
		#5;
		in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
		t0 = {3'd4, 3'd1, 3'd4, 3'd0, 3'd7, 3'd0, 3'd7, 3'd0, 3'd7, 3'd2, 3'd3, 3'd2, 3'd3, 3'd7, 3'd7, 3'd7};
		t1 = {3'd2, 3'd5, 3'd5, 3'd1, 3'd1, 3'd4, 3'd4, 3'd6, 3'd6, 3'd0, 3'd0, 3'd5, 3'd5, 3'd0, 3'd3, 3'd4};
		s0 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1};
		s1 = {1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0};
		//MAC result =  4290
		//-------------------------------
		#5;
		in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
		t0 = {3'd0, 3'd5, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0};
		t1 = {3'd0, 3'd0, 3'd5, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0};
		s0 = {1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
		s1 = {1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
		//MAC result =  961
		#5;
		in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
		t0 = {3'd0, 3'd3, 3'd4, 3'd7, 3'd0, 3'd3, 3'd4, 3'd7, 3'd0, 3'd3, 3'd4, 3'd7, 3'd1, 3'd3, 3'd1, 3'd3};
		t1 = {3'd0, 3'd0, 3'd0, 3'd0, 3'd2, 3'd2, 3'd2, 3'd2, 3'd4, 3'd4, 3'd4, 3'd4, 3'd0, 3'd0, 3'd3, 3'd3};
		s0 = {1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
		s1 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1};
		//MAC result =  -1379
		//-------------------------------
		#5;
		in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
		t0 = {3'd1, 3'd3, 3'd2, 3'd4, 3'd0, 3'd2, 3'd5, 3'd6, 3'd0, 3'd2, 3'd5, 3'd6, 3'd0, 3'd2, 3'd5, 3'd6};
		t1 = {3'd6, 3'd6, 3'd3, 3'd3, 3'd0, 3'd0, 3'd0, 3'd0, 3'd1, 3'd1, 3'd1, 3'd1, 3'd4, 3'd4, 3'd4, 3'd4};
		s0 = {1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
		s1 = {1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
		//MAC result =  1183
		//-------------------------------
		#5;
		in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
		t0 = {3'd1, 3'd3, 3'd4, 3'd7, 3'd1, 3'd3, 3'd4, 3'd7, 3'd0, 3'd7, 3'd0, 3'd7, 3'd0, 3'd7, 3'd2, 3'd3};
		t1 = {3'd0, 3'd0, 3'd0, 3'd0, 3'd7, 3'd7, 3'd7, 3'd7, 3'd1, 3'd1, 3'd4, 3'd4, 3'd6, 3'd6, 3'd0, 3'd0};
		s0 = {1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0};
		s1 = {1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1};
		//MAC result =  21324
		//-------------------------------
		#5;
		in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
		t0 = {3'd2, 3'd3, 3'd7, 3'd7, 3'd7, 3'd0, 3'd5, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0};
		t1 = {3'd5, 3'd5, 3'd0, 3'd3, 3'd4, 3'd0, 3'd0, 3'd5, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0};
		s0 = {1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
		s1 = {1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
		//MAC result =  -1599
		//-------------------------------
		#5;
		in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
		t0 = {3'd0, 3'd1, 3'd4, 3'd0, 3'd1, 3'd4, 3'd0, 3'd1, 3'd4, 3'd1, 3'd3, 3'd1, 3'd3, 3'd1, 3'd3, 3'd2};
		t1 = {3'd0, 3'd0, 3'd0, 3'd4, 3'd4, 3'd4, 3'd7, 3'd7, 3'd7, 3'd0, 3'd0, 3'd3, 3'd3, 3'd6, 3'd6, 3'd3};
		s0 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
		s1 = {1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0};
		//MAC result =  -2825
		//-------------------------------
		#5;
		in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
		t0 = {3'd4, 3'd0, 3'd0, 3'd0, 3'd1, 3'd4, 3'd1, 3'd4, 3'd2, 3'd4, 3'd2, 3'd4, 3'd2, 3'd4, 3'd0, 3'd3};
		t1 = {3'd3, 3'd0, 3'd1, 3'd4, 3'd2, 3'd2, 3'd3, 3'd3, 3'd1, 3'd1, 3'd4, 3'd4, 3'd6, 3'd6, 3'd0, 3'd0};
		s0 = {1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1};
		s1 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1};
		//MAC result =  282
		//-------------------------------
		#5;
		in_applied = {1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
		t0 = {3'd7, 3'd0, 3'd3, 3'd7, 3'd7, 3'd7, 3'd7, 3'd0, 3'd5, 3'd0, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0};
		t1 = {3'd0, 3'd5, 3'd5, 3'd5, 3'd0, 3'd3, 3'd4, 3'd0, 3'd0, 3'd5, 3'd5, 3'd0, 3'd0, 3'd0, 3'd0, 3'd0};
		s0 = {1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
		s1 = {1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1};
		//MAC result =  1761
		
    end
    
endmodule
